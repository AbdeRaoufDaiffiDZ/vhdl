library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity CLK_div is
generic(
period_max: integer := 50000000 -- max counting number for clock period
);
port(
clk: in std_logic; -- clock input;

clk_slow: out std_logic  -- clock output which gonna be slow when it will be devided

);
end CLK_div;


architecture arc of CLK_div is
signal clk_counter: integer:= 1;
signal tmp : std_logic := '0';

begin


divider: process(clk) 
	begin
	if(rising_edge(clk)) then
		clk_counter <= clk_counter + 1;

		if(clk_counter = period_max) then -- if the counter excied the max number return to 0
			tmp <= NOT tmp;
			clk_counter <= 1;

			
		end if;
		
	end if;
end  process;
clk_slow <= tmp;

end arc;